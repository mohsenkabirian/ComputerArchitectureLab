
module FuncTB;
reg a,b,c;
wire f;
func func_1(a,b,c,f);

////Making Clock
//initial
	//begin
	//	forever begin	
	//		clk=0;
	//		#10 clk = ~clk;
	//end
//end

endmodule
